-- #################################################################################################################################################################################
-- file :
--     gen_heartbeat.vhd
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- objective :
--     indicates FPGA activity.
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- level of description :
--     register tranfer level (RTL)
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- limitation :
--     clock ratio must be higher or equal to 16.
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- author :
--     Tugdual LE PELLETER
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- history :
--     2023-11-11
--         file creation
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- table of contents :
--     01. libraries
--     02. entity
--     03. architecture
--         03.01. constants
--         03.02. signals
--         03.03. input assignment
--         03.04. alive output pin generation
--         03.05. output assignment
-- #################################################################################################################################################################################

-- #################################################################################################################################################################################
-- 01. libraries
-- #################################################################################################################################################################################
    -- =============================================================================================================================================================================
	-- 01.01. standard
    -- =============================================================================================================================================================================
    library ieee;
        use ieee.std_logic_1164.all;
	    use ieee.numeric_std.all;
	    use ieee.math_real.all;

    -- =============================================================================================================================================================================
	-- 01.01. custom
    -- =============================================================================================================================================================================	
	library work;
	
-- #################################################################################################################################################################################
-- 02. entity
-- #################################################################################################################################################################################

entity ip_afifo_axis_top is
    port (
	     i_m_aclk    : in  std_logic
		;i_s_aclk    : in  std_logic
		;i_s_arst_n  : in  std_logic
		;i_s_data_en : in  std_logic
		;i_s_data    : in  std_logic_vector(7 downto 0)
		;o_m_data_en : out std_logic
		;o_m_data    : out std_logic_vector(7 downto 0)
		;o_ready     : out std_logic
	);
end entity ip_afifo_axis_top;

-- #################################################################################################################################################################################
-- 03. architecture
-- #################################################################################################################################################################################

architecture rtl of ip_afifo_axis_top is

    -- =============================================================================================================================================================================
	-- 03.01. components
    -- =============================================================================================================================================================================
    component ip_afifo_axis is
        port (
             wr_rst_busy   : out std_logic
            ;rd_rst_busy   : out std_logic
            ;m_aclk        : in  std_logic
            ;s_aclk        : in  std_logic
            ;s_aresetn     : in  std_logic
            ;s_axis_tvalid : in  std_logic
            ;s_axis_tready : out std_logic
            ;s_axis_tdata  : in  std_logic_vector(7 DOWNTO 0)
            ;s_axis_tuser  : in  std_logic_vector(3 DOWNTO 0)
            ;m_axis_tvalid : out std_logic
            ;m_axis_tready : in  std_logic
            ;m_axis_tdata  : out std_logic_vector(7 DOWNTO 0)
            ;m_axis_tuser  : out std_logic_vector(3 DOWNTO 0)
        );
    end component ip_afifo_axis;

    -- =============================================================================================================================================================================
	-- 03.01. constants
    -- =============================================================================================================================================================================

    -- =============================================================================================================================================================================
	-- 03.02. types
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.03. master (write)
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        type t_fsm_mst is (
	         state_fsm_mst_idle
		    ,state_fsm_mst_fifo_wr
	    );

    -- =============================================================================================================================================================================
	-- 03.02. signals
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.03. ip_afifo_axis
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        signal ip_afifo_axis_o_wr_rst_busy : std_logic;
        signal ip_afifo_axis_o_rd_rst_busy : std_logic;
        signal ip_afifo_axis_i_m_aclk      : std_logic;
        signal ip_afifo_axis_i_s_aclk      : std_logic;
        signal ip_afifo_axis_i_s_arst_n    : std_logic;
        signal ip_afifo_axis_i_s_tvalid    : std_logic;
        signal ip_afifo_axis_o_s_tready    : std_logic;
        signal ip_afifo_axis_i_s_tdata     : std_logic_vector(7 downto 0);
        signal ip_afifo_axis_i_s_tuser     : std_logic_vector(3 downto 0);
        signal ip_afifo_axis_o_m_tvalid    : std_logic;
        signal ip_afifo_axis_i_m_tready    : std_logic;
        signal ip_afifo_axis_o_m_tdata     : std_logic_vector(7 downto 0);
        signal ip_afifo_axis_o_m_tuser     : std_logic_vector(3 downto 0);
		signal s_fsm_fifo_wr               : t_fsm_mst;
		signal s_ready                     : std_logic;
		signal s_data                      : std_logic_vector(7 downto 0);
		signal s_data_en                   : std_logic;

begin

    -- =============================================================================================================================================================================
	-- 03.04. input assignment
    -- =============================================================================================================================================================================
    ip_afifo_axis_i_m_aclk   <= i_m_aclk;
    ip_afifo_axis_i_s_aclk   <= i_s_aclk;
    ip_afifo_axis_i_s_arst_n <= i_s_arst_n;
	s_data <= i_s_data;
	s_data_en <= i_s_data_en;

    -- =============================================================================================================================================================================
	-- 03.04. components
    -- =============================================================================================================================================================================
    inst_ip_afifo_axis : ip_afifo_axis
        port map (
             wr_rst_busy   => open
            ,rd_rst_busy   => open
            ,m_aclk        => ip_afifo_axis_i_m_aclk
            ,s_aclk        => ip_afifo_axis_i_s_aclk
            ,s_aresetn     => ip_afifo_axis_i_s_arst_n
            ,s_axis_tvalid => ip_afifo_axis_i_s_tvalid
            ,s_axis_tready => ip_afifo_axis_o_s_tready
            ,s_axis_tdata  => ip_afifo_axis_i_s_tdata
            ,s_axis_tuser  => ip_afifo_axis_i_s_tuser
            ,m_axis_tvalid => ip_afifo_axis_o_m_tvalid
            ,m_axis_tready => ip_afifo_axis_i_m_tready
            ,m_axis_tdata  => ip_afifo_axis_o_m_tdata
            ,m_axis_tuser  => ip_afifo_axis_o_m_tuser
        );

    -- =============================================================================================================================================================================
	-- 03.05. FSM FIFO write
    -- =============================================================================================================================================================================
    p_fsm_mst : process(ip_afifo_axis_i_m_aclk,ip_afifo_axis_i_s_arst_n)
	begin
	    if (ip_afifo_axis_i_s_arst_n = '0') then
		    s_fsm_fifo_wr <= state_fsm_mst_idle;
			s_ready <= '0';
			ip_afifo_axis_i_s_tdata <= (others => '0');
			ip_afifo_axis_i_s_tvalid <= '0';
			ip_afifo_axis_i_s_tuser <= (others => '0');
		elsif (rising_edge(ip_afifo_axis_i_m_aclk)) then
		    case s_fsm_fifo_wr is
			    when state_fsm_mst_idle =>
				    s_ready <= '1';
				    if (s_data_en = '1') then
					    s_fsm_fifo_wr <= state_fsm_mst_fifo_wr;
						s_ready <= '0';
						ip_afifo_axis_i_s_tdata <= s_data;
						--ip_afifo_axis_i_s_tvalid <= '1';
						ip_afifo_axis_i_s_tuser <= std_logic_vector(to_unsigned(4,ip_afifo_axis_i_s_tuser'length));
					end if;
				when state_fsm_mst_fifo_wr =>
				    -- wait for handshake
				    if (ip_afifo_axis_o_s_tready = '1') then
					    s_fsm_fifo_wr <= state_fsm_mst_idle;
					    ip_afifo_axis_i_s_tvalid <= '0';
						s_ready <= '1';
					end if;
			end case;
		end if;
	end process p_fsm_mst;

    -- =============================================================================================================================================================================
	-- 03.05. alive output pin generation
    -- =============================================================================================================================================================================

    -- =============================================================================================================================================================================
	-- 03.06. output assignment
    -- =============================================================================================================================================================================
    o_ready <= s_ready;
	ip_afifo_axis_i_m_tready <= '0';

end architecture rtl;

-- #################################################################################################################################################################################
-- EOF
-- #################################################################################################################################################################################