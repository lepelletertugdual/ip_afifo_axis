-- #################################################################################################################################################################################
-- file :
--     bch_ip_afifo_axis.vhd
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- objective :
--     gen_heartbeat.vhd testbench file.
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- level of description :
--     behavioral
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- limitation :
--     clock ratio must be higher or equal to 16.
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- author :
--     Tugdual LE PELLETER
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- history :
--     2023-11-11
--         file creation
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- table of contents :
--     01. libraries
--         01.01. standard
--         01.02. custom
--     02. entity
--     03. architecture
--         03.01. component declaration
--             03.01.01. DUT : gen_heartbeat
--         03.02. files
--             03.02.01. LOG
--             03.02.02. RPT
--         03.03. constants
--             03.03.01. SIM
--             03.03.02. DUT : gen_heartbeat
--             03.03.04. files
--         03.04. types
--             03.04.01. FSM
--                 03.04.01.01. fsm_main
--                 03.04.01.02. fsm_init
--                 03.04.01.03. fsm_test
--                 03.04.01.04. fsm_file_mgt_log
--                 03.04.01.05. fsm_file_mgt_rpt
--             03.04.02. test status
--         03.05. signals
--             03.05.01. SIM
--                 03.05.01.01. FSM
--                 03.05.01.02. files
--                 03.05.01.03. clock
--                 03.05.01.04. reset
--                 03.05.01.05. testbench
--             03.05.03. DUT : gen_heartbeat
--                 03.05.03.01. clock
--                 03.05.03.02. reset
--                 03.05.03.03. indicators
--         03.06. component instanciation
--             03.06.01. DUT : gen_heartbeat
--         03.07. reinit
--             03.07.01. SIM
--             03.07.02. DUT    
--         03.08. clock generation
--             03.08.01. DUT
--             03.08.02. SIM
--         03.09. fsm_main
--         03.10. fsm_init
--         03.11. fsm_test
--         03.12. fsm_file_mgt_log
--         03.13. fsm_file_mgt_rpt
--         03.14. simulation abort
-- #################################################################################################################################################################################

-- #################################################################################################################################################################################
-- 01. libraries
-- #################################################################################################################################################################################
    -- =============================================================================================================================================================================
	-- 01.01. standard
    -- =============================================================================================================================================================================
    library ieee;
        use ieee.std_logic_1164.all;
	    use ieee.numeric_std.all;
	    use ieee.math_real.all;
	
    library std;
        use std.textio.all;

    -- =============================================================================================================================================================================
	-- 01.02. custom
    -- =============================================================================================================================================================================
    library work;
        use work.pkg_mgt_file.all;
		use work.pkg_gen_heartbeat.all;
	
-- #################################################################################################################################################################################
-- 02. entity
-- #################################################################################################################################################################################

entity bch_ip_afifo_axis is
end entity bch_ip_afifo_axis;

-- #################################################################################################################################################################################
-- 03. architecture
-- #################################################################################################################################################################################

architecture behavioral of bch_ip_afifo_axis is

    -- =============================================================================================================================================================================
	-- 03.01. component declaration
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.01.01. DUT : gen_heartbeat
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        component gen_heartbeat is
            generic (
	             g_clk_i_freq : integer
		        ;g_clk_o_freq : integer
	        );
            port (
	             i_clk   : in  std_logic
		        ;i_rst   : in  std_logic
		        ;o_alive : out std_logic
				;o_error : out std_logic_vector(7 downto 0)
	        );
        end component gen_heartbeat;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.01.01. ip_afifo_axis
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
         component ip_afifo_axis is
             port (
                  wr_rst_busy   : out std_logic
                 ;rd_rst_busy   : out std_logic
                 ;m_aclk        : in  std_logic
                 ;s_aclk        : in  std_logic
                 ;s_aresetn     : in  std_logic
                 ;s_axis_tvalid : in  std_logic
                 ;s_axis_tready : out std_logic
                 ;s_axis_tdata  : in  std_logic_vector(7 DOWNTO 0)
                 ;s_axis_tuser  : in  std_logic_vector(3 DOWNTO 0)
                 ;m_axis_tvalid : out std_logic
                 ;m_axis_tready : in  std_logic
                 ;m_axis_tdata  : out std_logic_vector(7 DOWNTO 0)
                 ;m_axis_tuser  : out std_logic_vector(3 DOWNTO 0)
             );
         end component ip_afifo_axis;

    -- =============================================================================================================================================================================
	-- 03.02. files
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.02.01. LOG
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        file f_file_log : text;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.02.02. RPT
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        file f_file_rpt : text;

    -- =============================================================================================================================================================================
	-- 03.03. constants
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.01. SIM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    constant c_sim_clk_freq      : integer := 1_000_000_000;
	    constant c_sim_clk_delay     : time    := 0.9 us;
	    constant c_sim_rst_delay     : time    := 0.3 us;
        constant c_sim_clk_period_ns : time    := integer((real(1)/real(c_sim_clk_freq))*1.0e9)*1 ns;
	    constant c_sim_clk_period    : real    := real(1)/real(c_sim_clk_freq);
	
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.02. oscillator
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    constant c_osc_delay     : time := 2.4 us;
	    constant c_osc_freq      : integer := 100_000_000;
        constant c_osc_period_ns : time := integer((real(1)/real(c_osc_freq))*1.0e9)*1 ns;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.02. DUT : gen_heartbeat
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    constant c_dut_rst_delay    : time    := 2.5 us;
	    constant c_dut_clk_freq     : integer := c_osc_freq;
	    constant c_heartbeat_freq   : integer := 5_000_000;
		constant c_dut_clk_period   : real    := real(1)/real(c_dut_clk_freq);
	    constant c_heartbeat_period : real    := real(1)/real(c_heartbeat_freq);
	    constant c_alive_cycle_full : integer := integer(real(c_heartbeat_period)/real(c_sim_clk_period));
	    constant c_alive_cycle_half : integer := integer(real(c_alive_cycle_full)/real(2));
	
		-- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.02. ip_afifo_axis
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    constant c_ip_fifo_arst_n_delay      : time    := 1.2 us;
		constant c_ip_fifo_depth             : integer := 128;
		constant c_ip_fifo_data_width        : integer := 8;
		constant c_ip_fifo_clk_freq_wr       : integer := 1_000_000;
		constant c_ip_fifo_clk_freq_wr_delay : time    := 0.3 us;
		constant c_ip_fifo_clk_freq_rd       : integer := 1_000_000;
		constant c_ip_fifo_clk_freq_rd_delay : time    := 1.0 us;
		constant c_ip_fifo_period_wr_ns      : time    := integer((real(1)/real(c_ip_fifo_clk_freq_wr))*1.0e9)*1 ns;
		constant c_ip_fifo_period_rd_ns      : time    := integer((real(1)/real(c_ip_fifo_clk_freq_rd))*1.0e9)*1 ns;
		constant c_ratio_clk_sim_clk_wr      : integer := integer(real(c_sim_clk_freq)/real(c_ip_fifo_clk_freq_wr));
		constant c_ratio_clk_sim_clk_rd      : integer := integer(real(c_sim_clk_freq)/real(c_ip_fifo_clk_freq_rd));
	
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.03. simulation duration
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		constant c_sim_duration_factor : integer := 16;
	    constant c_sim_duration_ns     : integer := integer(real(c_sim_duration_factor)*real(c_heartbeat_period)/real(c_sim_clk_period));
	
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.04. file
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		constant c_file_log_name : string := "log_bch_ip_afifo_axis_wrapper_nexys_a7_sim.csv";
		constant c_file_rpt_name : string := "rpt_bch_ip_afifo_axis_wrapper_nexys_a7_sim.txt";
	
    -- =============================================================================================================================================================================
	-- 03.04. types
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.01. FSM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		    -- =====================================================================================================================================================================
			-- 03.04.01.01. fsm_main
			-- =====================================================================================================================================================================
	        type t_fsm_main is (
	             state_fsm_main_start
                ,state_fsm_main_file_rpt_open
                ,state_fsm_main_file_log_open
			    ,state_fsm_main_init
		        ,state_fsm_main_run
                ,state_fsm_main_file_rpt_close
                ,state_fsm_main_file_log_close
		        ,state_fsm_main_stop
	        );

		    -- =====================================================================================================================================================================
			-- 03.04.01.02. fsm_init
			-- =====================================================================================================================================================================
	        type t_fsm_init is (
	             state_fsm_init_idle
		        ,state_fsm_init_run
		        ,state_fsm_init_done
	        );

		    -- =====================================================================================================================================================================
			-- 03.04.01.03. fsm_test
			-- =====================================================================================================================================================================
	        type t_fsm_test is (
	             state_fsm_test_idle
				,state_fsm_test_run_fifo_wr
				,state_fsm_test_run_fifo_rd
				,state_fsm_test_run_check
		        ,state_fsm_test_done
	        );

		    -- =====================================================================================================================================================================
			-- 03.04.01.03. fsm_test_fifo_wr
			-- =====================================================================================================================================================================
	        type t_fsm_test_fifo_wr is (
	             state_fsm_test_run_fifo_idle
				,state_fsm_test_run_fifo_wr
		        ,state_fsm_test_run_fifo_done
	        );

		    -- =====================================================================================================================================================================
			-- 03.04.01.03. fsm_test_fifo_rd
			-- =====================================================================================================================================================================
	        type t_fsm_test_fifo_rd is (
	             state_fsm_test_run_fifo_idle
				,state_fsm_test_run_fifo_rd
		        ,state_fsm_test_run_fifo_done
	        );
	
		    -- =====================================================================================================================================================================
			-- 03.04.01.04. fsm_file_mgt_log
			-- =====================================================================================================================================================================
	        type t_fsm_file_mgt_log is (
	             state_fsm_file_mgt_log_open
				,state_fsm_file_mgt_log_write_head
	            ,state_fsm_file_mgt_log_write_data
		        ,state_fsm_file_mgt_log_close
				,state_fsm_file_mgt_log_done
	        );

		    -- =====================================================================================================================================================================
			-- 03.04.01.04. fsm_file_mgt_rpt
			-- =====================================================================================================================================================================
	        type t_fsm_file_mgt_rpt is (
	             state_fsm_file_mgt_rpt_open
	            ,state_fsm_file_mgt_rpt_write_status
		        ,state_fsm_file_mgt_rpt_close
				,state_fsm_file_mgt_rpt_done
	        );

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.02. test status
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	        type t_sim_test_status is (
	             TEST_OK
	            ,TEST_KO
	        );

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.01. Arrays
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        type t_array is array (integer range <>) of std_logic_vector(c_ip_fifo_data_width-1 downto 0);
	
    -- =============================================================================================================================================================================
	-- 03.05. signals
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.02. SIM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		    -- =====================================================================================================================================================================
			-- 03.05.02.01. FSM
			-- =====================================================================================================================================================================
	        signal s_fsm_main_state   : t_fsm_main;
	        signal s_fsm_init_state   : t_fsm_init;
	        signal s_fsm_test_state   : t_fsm_test;
			signal s_fsm_test_fifo_wr_state : t_fsm_test_fifo_wr;
			signal s_fsm_test_fifo_rd_state : t_fsm_test_fifo_rd;
		    signal s_fsm_file_mgt_log : t_fsm_file_mgt_log;
		    signal s_fsm_file_mgt_rpt : t_fsm_file_mgt_rpt;
	
		    -- =====================================================================================================================================================================
			-- 03.05.02.02. files
			-- =====================================================================================================================================================================
		    signal s_sim_file_req_log_open  : std_logic;
		    signal s_sim_file_ack_log_open  : std_logic;
		    signal s_sim_file_req_log_close : std_logic;
		    signal s_sim_file_ack_log_close : std_logic;
		    signal s_sim_file_req_rpt_open  : std_logic;
		    signal s_sim_file_ack_rpt_open  : std_logic;
		    signal s_sim_file_req_rpt_close : std_logic;
		    signal s_sim_file_ack_rpt_close : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.02.03. clock
			-- =====================================================================================================================================================================
            signal s_sim_clk : std_logic;
	        signal s_osc     : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.02.04. reset
			-- =====================================================================================================================================================================
		    signal s_sim_rst : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.02.05. testbench
			-- =====================================================================================================================================================================
	        signal s_sim_cnt         : integer range 0 to c_sim_duration_ns-1;
		    signal s_sim_done        : std_logic;
		    signal s_sim_init_req    : std_logic;
		    signal s_sim_init_ack    : std_logic;
		    signal s_sim_test_req    : std_logic;
		    signal s_sim_test_ack    : std_logic;
			signal s_sim_test_fifo_wr_req : std_logic;
			signal s_sim_test_fifo_wr_ack : std_logic;
			signal s_sim_test_fifo_wr_req_reg : std_logic_vector(c_ratio_clk_sim_clk_wr-1 downto 0);
			signal s_sim_test_fifo_wr_req_reg_gen_tmp : std_logic_vector(c_ratio_clk_sim_clk_wr-1 downto 0);
			signal s_sim_test_fifo_wr_req_reg_gen : std_logic;
			signal s_sim_test_fifo_rd_req : std_logic;
			signal s_sim_test_fifo_rd_ack : std_logic;
			signal s_sim_test_fifo_rd_req_reg : std_logic_vector(c_ratio_clk_sim_clk_rd-1 downto 0);
			signal s_sim_test_fifo_rd_req_reg_gen_tmp : std_logic_vector(c_ratio_clk_sim_clk_rd-1 downto 0);
			signal s_sim_test_fifo_rd_req_reg_gen : std_logic;
		    signal s_sim_test_status : t_sim_test_status;
			signal s_error           : std_logic;
			signal s_array_data      : t_array(0 to c_ip_fifo_depth-1);
			signal s_array_data_rd      : t_array(0 to c_ip_fifo_depth-1);
			signal s_array_data_idx  : integer range 0 to c_ip_fifo_depth-1;
			signal s_array_data_cnt  : integer range 0 to c_ip_fifo_depth-1;
			signal s_ip_fifo_axis_clk_wr : std_logic;
			signal s_ip_fifo_axis_clk_rd : std_logic;
			signal s_ip_afifo_axis_data_idx_wr : integer range 0 to c_ip_fifo_depth-1;
			signal s_ip_afifo_axis_data_idx_rd : integer range 0 to c_ip_fifo_depth-1;
			signal s_ip_afifo_axis_data_idx_check : integer range 0 to c_ip_fifo_depth-1;
			signal s_error_data_check : std_logic;
	
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.03. DUT : gen_heartbeat
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        signal s_dut_i_clk   : std_logic;
	    signal s_dut_i_rst   : std_logic;
		signal s_dut_o_alive : std_logic;
		signal s_dut_o_error : std_logic_vector(7 downto 0);

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.03. ip_afifo_axis
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        signal s_ip_afifo_axis_i_m_aclk   : std_logic; -- write
        signal s_ip_afifo_axis_i_s_aclk   : std_logic; -- read
        signal s_ip_afifo_axis_i_s_arst_n : std_logic;
        signal s_ip_afifo_axis_i_s_tvalid : std_logic;
        signal s_ip_afifo_axis_o_s_tready : std_logic;
        signal s_ip_afifo_axis_i_s_tdata  : std_logic_vector(7 downto 0);
        signal s_ip_afifo_axis_i_s_tuser  : std_logic_vector(3 downto 0);
        signal s_ip_afifo_axis_o_m_tvalid : std_logic;
        signal s_ip_afifo_axis_i_m_tready : std_logic;
        signal s_ip_afifo_axis_o_m_tdata  : std_logic_vector(7 downto 0);
        signal s_ip_afifo_axis_o_m_tuser  : std_logic_vector(3 downto 0);

begin

    -- =============================================================================================================================================================================
	-- 03.07. reset management
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.07.01. SIM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_sim_rst <= '1','0' after c_sim_rst_delay;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.07.02. DUT
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_dut_i_rst <= '1','0' after c_dut_rst_delay;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.07.02. ip_afifo_axis
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_ip_afifo_axis_i_s_arst_n <= '0','1' after c_ip_fifo_arst_n_delay;

    -- =============================================================================================================================================================================
	-- 03.08. clock generation
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.08.01. SIM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    p_gen_sim_clk : process
		begin
	        s_sim_clk <= '0';
	        wait for c_sim_clk_delay;
		    while true loop
		        s_sim_clk <= '1';
			    wait for c_sim_clk_period_ns/2;
			    s_sim_clk <= '0';
			    wait for c_sim_clk_period_ns/2;
		    end loop;
	    end process p_gen_sim_clk;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.08.02. oscillator
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    p_gen_osc : process
		begin
	        s_osc <= '0';
	        wait for c_osc_delay;
		    while true loop
		        s_osc <= '1';
			    wait for c_osc_period_ns/2;
			    s_osc <= '0';
			    wait for c_osc_period_ns/2;
		    end loop;
	    end process p_gen_osc;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.08.02. ip_fifo_axis write clock (slave)
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    p_gen_ip_afifo_axis_wr_clk : process
		begin
	        s_ip_fifo_axis_clk_wr <= '0';
	        wait for c_ip_fifo_clk_freq_wr_delay;
		    while true loop
		        s_ip_fifo_axis_clk_wr <= '1';
			    wait for c_ip_fifo_period_wr_ns/2;
			    s_ip_fifo_axis_clk_wr <= '0';
			    wait for c_ip_fifo_period_wr_ns/2;
		    end loop;
	    end process p_gen_ip_afifo_axis_wr_clk;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.08.02. ip_fifo_axis read clock (master)
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    p_gen_ip_afifo_axis_rd_clk : process
		begin
	        s_ip_fifo_axis_clk_rd <= '0';
	        wait for c_ip_fifo_clk_freq_rd_delay;
		    while true loop
		        s_ip_fifo_axis_clk_rd <= '1';
			    wait for c_ip_fifo_period_rd_ns/2;
			    s_ip_fifo_axis_clk_rd <= '0';
			    wait for c_ip_fifo_period_rd_ns/2;
		    end loop;
	    end process p_gen_ip_afifo_axis_rd_clk;

    -- =============================================================================================================================================================================
	-- 03.08. clock assignment
    -- =============================================================================================================================================================================
    s_dut_i_clk <= s_osc;
	s_ip_afifo_axis_i_s_aclk <= s_ip_fifo_axis_clk_wr;
	s_ip_afifo_axis_i_m_aclk <= s_ip_fifo_axis_clk_rd;

    -- =============================================================================================================================================================================
	-- 03.06. component instanciation
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.06.02. DUT : gen_heartbeat
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        inst_dut_gen_heartbeat : gen_heartbeat
            generic map (
	             g_clk_i_freq => c_dut_clk_freq
		        ,g_clk_o_freq => c_heartbeat_freq
	        )
            port map (
	             i_clk   => s_dut_i_clk
		        ,i_rst   => s_dut_i_rst
		        ,o_alive => s_dut_o_alive
				,o_error => s_dut_o_error
	        );
			
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.01.01. ip_afifo_axis
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        inst_ip_afifo_axis : ip_afifo_axis
            port map (
                 wr_rst_busy   => open
                ,rd_rst_busy   => open
                ,m_aclk        => s_ip_afifo_axis_i_m_aclk
                ,s_aclk        => s_ip_afifo_axis_i_s_aclk
                ,s_aresetn     => s_ip_afifo_axis_i_s_arst_n
                ,s_axis_tvalid => s_ip_afifo_axis_i_s_tvalid
                ,s_axis_tready => s_ip_afifo_axis_o_s_tready
                ,s_axis_tdata  => s_ip_afifo_axis_i_s_tdata
                ,s_axis_tuser  => s_ip_afifo_axis_i_s_tuser
                ,m_axis_tvalid => s_ip_afifo_axis_o_m_tvalid
                ,m_axis_tready => s_ip_afifo_axis_i_m_tready
                ,m_axis_tdata  => s_ip_afifo_axis_o_m_tdata
                ,m_axis_tuser  => s_ip_afifo_axis_o_m_tuser
            );
	     		
    -- =============================================================================================================================================================================
	-- 03.09. fsm_main
    -- =============================================================================================================================================================================
	p_fsm_main : process(s_sim_rst,s_sim_clk)
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_main_state <= state_fsm_main_start;
			s_sim_done <= '0';
			s_sim_init_req <= '0';
			s_sim_test_req <= '0';
			s_sim_file_req_log_open <= '0';
			s_sim_file_req_log_close <= '0';
			s_sim_file_req_rpt_open <= '0';
			s_sim_file_req_rpt_close <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_done <= '0';
            s_sim_init_req <= '0';
			s_sim_test_req <= '0';
			s_sim_file_req_log_open <= '0';
			s_sim_file_req_log_close <= '0';
			s_sim_file_req_rpt_open <= '0';
			s_sim_file_req_rpt_close <= '0';
		    case s_fsm_main_state is
			    -- wait for DUT reset deassertion
				when state_fsm_main_start =>
				    if (s_dut_i_rst = '0') then
					    s_fsm_main_state <= state_fsm_main_file_rpt_open;
						s_sim_file_req_rpt_open <= '1';
					end if;
				-- wait for RPT file to be opened
			    when state_fsm_main_file_rpt_open =>
				    if (s_sim_file_ack_rpt_open = '1') then
					    s_fsm_main_state <= state_fsm_main_file_log_open;
					    s_sim_file_req_log_open <= '1';
					end if;
				-- wait for LOG file to be opened
				when state_fsm_main_file_log_open =>
				    if (s_sim_file_ack_log_open = '1') then
					    s_fsm_main_state <= state_fsm_main_init;
						s_sim_init_req <= '1';
					end if;
				-- waiting for init done
				when state_fsm_main_init =>
				    if (s_sim_init_ack = '1') then
					    s_fsm_main_state <= state_fsm_main_run;
					    s_sim_test_req <= '1';
					end if;
				-- waiting for test done
				when state_fsm_main_run =>
                    if (s_sim_test_ack = '1') then
					    s_fsm_main_state <= state_fsm_main_file_log_close;
						s_sim_file_req_log_close <= '1';
					end if;
				-- waiting for data file to be closed
				when state_fsm_main_file_log_close =>
                    if (s_sim_file_ack_log_close = '1') then
					    s_fsm_main_state <= state_fsm_main_file_rpt_close;
						s_sim_file_req_rpt_close <= '1';
					end if;
				-- waiting for SIM report file to be closed
				when state_fsm_main_file_rpt_close =>
                    if (s_sim_file_ack_rpt_close = '1') then
					    s_fsm_main_state <= state_fsm_main_stop;
				        s_sim_done <= '1';
					end if;
				-- test stopped
                when state_fsm_main_stop =>
                    null;
			end case;
		end if;
	end process p_fsm_main;

    -- =============================================================================================================================================================================
	-- 03.10. fsm_init
    -- =============================================================================================================================================================================
	fsm_init : process(s_sim_rst,s_sim_clk)
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_init_state <= state_fsm_init_idle;
			s_sim_init_ack <= '0';
			s_array_data_cnt <= 0;
			s_array_data_idx <= 0;
			s_array_data <= (others => (others => '0'));
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_init_ack <= '0';
		    case s_fsm_init_state is
			    -- waiting for init request
			    when state_fsm_init_idle =>
				    if (s_sim_init_req = '1') then
					    s_fsm_init_state <= state_fsm_init_run;
					end if;
				-- running init
				when state_fsm_init_run =>
					s_array_data(s_array_data_idx) <= std_logic_vector(to_unsigned(s_array_data_cnt,c_ip_fifo_data_width));
					if (s_array_data_idx = c_ip_fifo_depth-1) then
					    s_array_data_idx <= 0;
						s_array_data_cnt <= 0;
					    s_fsm_init_state <= state_fsm_init_done;
                        s_sim_init_ack <= '1';
					else
						s_array_data_cnt <= s_array_data_cnt + 1;
					    s_array_data_idx <= s_array_data_idx + 1;
					end if;
				-- init done
                when state_fsm_init_done =>
				    null;
			end case;
		end if;
	end process fsm_init;

    -- =============================================================================================================================================================================
	-- 03.11. fsm_test
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.06.02. main
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    p_fsm_test_main : process(s_sim_rst,s_sim_clk)
	    begin
	        if (s_sim_rst = '1') then
	    	    s_fsm_test_state <= state_fsm_test_idle;
	    		s_sim_cnt <= 0;
	    		s_sim_test_ack <= '0';
	    		s_sim_test_status <= TEST_OK;
	    		s_sim_test_fifo_wr_req <= '0';
                s_sim_test_fifo_rd_req <= '0';
				s_ip_afifo_axis_data_idx_check <= 0;
				s_error_data_check <= '0';
	    	elsif (rising_edge(s_sim_clk)) then
	    	    s_sim_test_ack <= '0';
	    		s_sim_test_fifo_wr_req <= '0';
                s_sim_test_fifo_rd_req <= '0';
	    	    case s_fsm_test_state is
	    		    -- waiting for test request
	    		    when state_fsm_test_idle =>
	    			    if (s_sim_test_req = '1') then
	    				    s_fsm_test_state <= state_fsm_test_run_fifo_wr;
	    					s_sim_test_fifo_wr_req <= '1';
	    				end if;
	    			-- running test
	    			when state_fsm_test_run_fifo_wr =>
	    			    if (s_sim_test_fifo_wr_ack = '1') then
	    				    s_fsm_test_state <= state_fsm_test_run_fifo_rd;
							s_sim_test_fifo_rd_req <= '1';
						end if;
	    			when state_fsm_test_run_fifo_rd =>
	    			    if (s_sim_test_fifo_rd_ack = '1') then
						    s_fsm_test_state <= state_fsm_test_run_check;
						end if;
					when state_fsm_test_run_check =>
					    -- verification
					    if (s_array_data(s_ip_afifo_axis_data_idx_check) /= s_array_data_rd(s_ip_afifo_axis_data_idx_check)) then
						    s_error_data_check <= '1';
						end if;
						-- index incrementation
					    if (s_ip_afifo_axis_data_idx_check = c_ip_fifo_depth-1) then
						    s_fsm_test_state <= state_fsm_test_done;
							s_sim_test_ack <= '1';
						    s_ip_afifo_axis_data_idx_check <= 0;
							if (s_error_data_check = '0') then
							    s_sim_test_status <= TEST_OK;
							else
							    s_sim_test_status <= TEST_KO;
							end if;
						else
						    s_ip_afifo_axis_data_idx_check <= s_ip_afifo_axis_data_idx_check + 1;
						end if;
                    when state_fsm_test_done =>
                        null;
	    		end case;
	    	end if;
	    end process p_fsm_test_main;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.06.02. write asynchronous FIFO 
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        p_fifo_wr_req_sr: process(s_sim_rst,s_sim_clk)
		begin
		    if (s_sim_rst = '1') then
			    s_sim_test_fifo_wr_req_reg <= (others => '0');
			elsif (rising_edge(s_sim_clk)) then
			    s_sim_test_fifo_wr_req_reg <= s_sim_test_fifo_wr_req_reg(s_sim_test_fifo_wr_req_reg'length-2 downto 0) & s_sim_test_fifo_wr_req;
			end if;
		end process p_fifo_wr_req_sr;
 
        s_sim_test_fifo_wr_req_reg_gen_tmp(0) <= s_sim_test_fifo_wr_req_reg(0);
		or_gen_wr_req : for i in 1 to c_ratio_clk_sim_clk_wr-1 generate
		    s_sim_test_fifo_wr_req_reg_gen_tmp(i) <= s_sim_test_fifo_wr_req_reg(i) or s_sim_test_fifo_wr_req_reg_gen_tmp(i-1);
		end generate or_gen_wr_req;
		s_sim_test_fifo_wr_req_reg_gen <= s_sim_test_fifo_wr_req_reg_gen_tmp(s_sim_test_fifo_wr_req_reg_gen_tmp'length-1);
 
        p_fsm_test_run_fifo_wr : process(s_ip_fifo_axis_clk_wr,s_ip_afifo_axis_i_s_arst_n)
		begin
		    if (s_ip_afifo_axis_i_s_arst_n = '0') then
			    s_fsm_test_fifo_wr_state <= state_fsm_test_run_fifo_idle;
				s_ip_afifo_axis_i_s_tdata <= (others => '0');
                s_ip_afifo_axis_i_s_tvalid <= '0';
				s_ip_afifo_axis_data_idx_wr <= 0;
				s_ip_afifo_axis_i_s_tuser <= (others => '0');
				s_sim_test_fifo_wr_ack <= '0';
			elsif (rising_edge(s_ip_fifo_axis_clk_wr)) then
				s_ip_afifo_axis_i_s_tvalid <= '0';
				s_sim_test_fifo_wr_ack <= '0';
			    case s_fsm_test_fifo_wr_state is
				    when state_fsm_test_run_fifo_idle =>
					    if (s_sim_test_fifo_wr_req_reg_gen = '1') then
					        s_fsm_test_fifo_wr_state <= state_fsm_test_run_fifo_wr;
						end if;
					when state_fsm_test_run_fifo_wr =>
					    if (s_ip_afifo_axis_o_s_tready = '1') then
						    -- handshake
						    s_ip_afifo_axis_i_s_tvalid <= '1';
					        s_ip_afifo_axis_i_s_tdata <= s_array_data(s_ip_afifo_axis_data_idx_wr);
					        if (s_ip_afifo_axis_data_idx_wr = c_ip_fifo_depth-1) then
					            s_fsm_test_fifo_wr_state <= state_fsm_test_run_fifo_done;
								s_ip_afifo_axis_data_idx_wr <= 0;
								s_sim_test_fifo_wr_ack <= '1';
					        else
					            s_ip_afifo_axis_data_idx_wr <= s_ip_afifo_axis_data_idx_wr + 1;
					        end if;
					    end if;
					 when state_fsm_test_run_fifo_done =>
					     null;
				end case;
			end if;
		end process p_fsm_test_run_fifo_wr;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.06.02. read asynchronous FIFO 
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        p_fifo_rd_req_sr: process(s_sim_rst,s_sim_clk)
		begin
		    if (s_sim_rst = '1') then
			     s_sim_test_fifo_rd_req_reg <= (others => '0');
			elsif (rising_edge(s_sim_clk)) then
			    s_sim_test_fifo_rd_req_reg <= s_sim_test_fifo_rd_req_reg(s_sim_test_fifo_rd_req_reg'length-2 downto 0) & s_sim_test_fifo_rd_req;
			end if;
		end process p_fifo_rd_req_sr;
 
        s_sim_test_fifo_rd_req_reg_gen_tmp(0) <= s_sim_test_fifo_rd_req_reg(0);
		or_gen_rd_req : for i in 1 to c_ratio_clk_sim_clk_rd-1 generate
		    s_sim_test_fifo_rd_req_reg_gen_tmp(i) <= s_sim_test_fifo_rd_req_reg(i) or s_sim_test_fifo_rd_req_reg_gen_tmp(i-1);
		end generate or_gen_rd_req;
		s_sim_test_fifo_rd_req_reg_gen <= s_sim_test_fifo_rd_req_reg_gen_tmp(s_sim_test_fifo_rd_req_reg_gen_tmp'length-1);
 
        p_fsm_test_run_fifo_rd : process(s_ip_fifo_axis_clk_rd,s_ip_afifo_axis_i_s_arst_n)
		begin
		    if (s_ip_afifo_axis_i_s_arst_n = '0') then
			    s_fsm_test_fifo_rd_state <= state_fsm_test_run_fifo_idle;
				s_ip_afifo_axis_data_idx_rd <= 0;
				s_ip_afifo_axis_i_m_tready <= '0';
				s_array_data_rd <= (others => (others => '0'));
				s_sim_test_fifo_rd_ack <= '0';
			elsif (rising_edge(s_ip_fifo_axis_clk_rd)) then
				s_sim_test_fifo_rd_ack <= '0';
			    case s_fsm_test_fifo_rd_state is
				    when state_fsm_test_run_fifo_idle =>
					    if (s_sim_test_fifo_rd_req_reg_gen = '1') then
					        s_fsm_test_fifo_rd_state <= state_fsm_test_run_fifo_rd;
							-- anticipating read latency (1 clock period)
				            s_ip_afifo_axis_i_m_tready <= '1';
						end if;
					when state_fsm_test_run_fifo_rd =>
						-- handshake
					    if (s_ip_afifo_axis_o_m_tvalid = '1') then
					        s_array_data_rd(s_ip_afifo_axis_data_idx_rd) <= s_ip_afifo_axis_o_m_tdata;
					        if (s_ip_afifo_axis_data_idx_rd = c_ip_fifo_depth-1) then
					            s_fsm_test_fifo_rd_state <= state_fsm_test_run_fifo_done;
								s_ip_afifo_axis_data_idx_rd <= 0;
								s_sim_test_fifo_rd_ack <= '1';
				                s_ip_afifo_axis_i_m_tready <= '0';
					        else
					            s_ip_afifo_axis_data_idx_rd <= s_ip_afifo_axis_data_idx_rd + 1;
					        end if;
					    end if;
					 when state_fsm_test_run_fifo_done =>
					     null;
				end case;
			end if;
		end process p_fsm_test_run_fifo_rd;

    -- =============================================================================================================================================================================
	-- 03.12. fsm_file_mgt_log
    -- =============================================================================================================================================================================
	p_fsm_file_mgt_log : process(s_sim_rst,s_sim_clk)
		constant c_justified  : side   := right;
		constant c_field      : width  := 0;
		constant c_unit       : time   := ns;
		constant c_separator  : string := ",";
		constant c_value_head : string := "time,data";
	    variable v_value_time : time;
		variable v_value_data : string(1 to 4);
		variable v_value_foot : string(1 to 7);
		variable v_line       : line;
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_open;
		    s_sim_file_ack_log_open <= '0';
			s_sim_file_ack_log_close <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_file_ack_log_open <= '0';
			s_sim_file_ack_log_close <= '0';
            case s_fsm_file_mgt_log is
                -- open file
			    when state_fsm_file_mgt_log_open =>
				    if (s_sim_file_req_log_open = '1') then
					    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_write_head;
						s_sim_file_ack_log_open <= '1';
						proc_file_log_open(c_file_log_name,f_file_log);
					end if;
				-- write header
				when state_fsm_file_mgt_log_write_head =>
					    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_write_data;
						write(v_line,c_value_head,c_justified,c_field);
	                    writeline(f_file_log,v_line);
				-- write data
				when state_fsm_file_mgt_log_write_data =>
				    if (s_sim_file_req_log_close = '1') then
					    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_close;
						-- timestamp
						v_value_time := now;
						write(v_line,v_value_time,c_justified,c_field,c_unit);
						-- separator
						write(v_line,c_separator,c_justified,c_field);
						-- data value
						v_value_data := "NONE";
					    write(v_line,v_value_data,c_justified,c_field);
	                    writeline(f_file_log,v_line);
					end if;
                -- close file
				when state_fsm_file_mgt_log_close =>
					s_fsm_file_mgt_log <= state_fsm_file_mgt_log_done;
				    s_sim_file_ack_log_close <= '1';
                    proc_file_log_close(c_file_log_name,f_file_log);
				-- done
				when state_fsm_file_mgt_log_done  =>
				    null;
			end case;
		end if;
	end process p_fsm_file_mgt_log;

    -- =============================================================================================================================================================================
	-- 03.13. fsm_file_mgt_rpt
    -- =============================================================================================================================================================================
	p_fsm_file_mgt_rpt : process(s_sim_rst,s_sim_clk)
		constant c_justified    : side  := right;
		constant c_field        : width := 0;
		variable v_value_status : string(1 to 7);
		variable v_line         : line;
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_open;
		    s_sim_file_ack_rpt_open <= '0';
			s_sim_file_ack_rpt_close <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_file_ack_rpt_open <= '0';
			s_sim_file_ack_rpt_close <= '0';
            case s_fsm_file_mgt_rpt is
                -- open file
			    when state_fsm_file_mgt_rpt_open =>
				    if (s_sim_file_req_rpt_open = '1') then
					    s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_write_status;
						s_sim_file_ack_rpt_open <= '1';
						proc_file_rpt_open(c_file_rpt_name,f_file_rpt);
					end if;
				-- write status
				when state_fsm_file_mgt_rpt_write_status =>
				    if (s_sim_file_req_rpt_close = '1') then
					    s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_close;
					    -- write test status
					    case s_sim_test_status is
					        when TEST_OK => v_value_status := "TEST_OK";
						    when others  => v_value_status := "TEST_KO";
					    end case;
					    write(v_line,v_value_status,c_justified,c_field);
	                    writeline(f_file_rpt,v_line);
					end if;
                -- close file
				when state_fsm_file_mgt_rpt_close =>
					s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_done;
				    s_sim_file_ack_rpt_close <= '1';
                    proc_file_rpt_close(c_file_rpt_name,f_file_rpt);
				-- done
				when state_fsm_file_mgt_rpt_done  =>
				    null;
			end case;
		end if;
	end process p_fsm_file_mgt_rpt;

    -- =============================================================================================================================================================================
	-- 03.14. error detection
    -- =============================================================================================================================================================================
	p_check_dut_error : process(s_dut_i_rst,s_sim_clk)
	    variable v_error : std_logic;
	begin
	    if (s_dut_i_rst = '1') then
	        v_error := '0';
			s_error <= '0';
	    elsif (rising_edge(s_sim_clk)) then
		    v_error := '0';
			-- parsing error vector
		    for i in 0 to s_dut_o_error'length-1 loop
		        -- error detected
			    if (s_dut_o_error(i) = '1') then
				    v_error := '1';
				end if;
			end loop;
			s_error <= v_error;
		end if;
	end process p_check_dut_error;	
	
    -- =============================================================================================================================================================================
	-- 03.14. simulation abort : clock ratio error
    -- =============================================================================================================================================================================
	p_sim_abort : process(s_sim_clk)
	begin
		if (rising_edge(s_sim_clk)) then
            if (s_error = '1') then
			    assert false 
				    report "end of simulation - DUT error detected" 
					    severity failure;
			end if;
			if (s_error_data_check = '1') then
			    assert false 
				    report "end of simulation - data arrays are not identical" 
					    severity failure;
			end if;
		end if;
	end process p_sim_abort;

    -- =============================================================================================================================================================================
	-- 03.14. end of simulation
    -- =============================================================================================================================================================================
	p_sim_end : process(s_sim_clk)
	begin
		if (rising_edge(s_sim_clk)) then
            if (s_sim_done = '1') then
			    assert false 
				    report "end of simulation - success" 
					    severity failure;
			end if;
		end if;
	end process p_sim_end;

end architecture behavioral;

-- #################################################################################################################################################################################
-- EOF
-- #################################################################################################################################################################################